module alu #(
    parameter WIDTH = 16
)(
    input  logic     ALUop1,      // clock 
    input  logic     ALUop2,      // reset
    input  logic     ALUctrl,
    output logic     SUM,
    output logic     EQ  // output
);



endmodule
