module top#(
    parameter ADDRESS_WIDTH = 32,
    DATA_WIDTH = 32
)(

);



topAlu alu(

);

pctop myPC(

);