module controlunit(
    input logic [2:0]   funct3_i,
    input logic         funct7_i,
    input logic [6:0]   op_i,
    output logic        mem_write,
    output logic        alu_src,
    

    

)