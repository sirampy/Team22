// reg from Exectute to store in memory

module regEtoS #(
        parameter ADDRESS_WIDTH = 32,
              DATA_WIDTH = 32
)(
    input logic clk_i,
    //control inputs

    //other inputs

    //control outputs

    //other outputs
);