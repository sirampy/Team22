module top#(
    parameter ADDRESS_WIDTH = ,
    DATA_WIDTH = 
)(

);



topAlu alu(

);

pctop myPC(

);