module top#(
    parameter ADDRESS_WIDTH = 32,
    DATA_WIDTH = 32
)(

);



topAku alu(

);

pctop myPC(

);